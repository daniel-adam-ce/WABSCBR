// DE2_115_Qsys.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module DE2_115_Qsys (
		input  wire [3:0]  button_pio_external_connection_export, // button_pio_external_connection.export
		input  wire        clk_100_clk_in_clk,                    //                 clk_100_clk_in.clk
		input  wire        clk_100_clk_in_reset_reset_n,          //           clk_100_clk_in_reset.reset_n
		input  wire        clk_io_clk_in_clk,                     //                  clk_io_clk_in.clk
		inout  wire [15:0] cy7c67200_if_0_conduit_end_DATA,       //     cy7c67200_if_0_conduit_end.DATA
		output wire [1:0]  cy7c67200_if_0_conduit_end_ADDR,       //                               .ADDR
		output wire        cy7c67200_if_0_conduit_end_RD_N,       //                               .RD_N
		output wire        cy7c67200_if_0_conduit_end_WR_N,       //                               .WR_N
		output wire        cy7c67200_if_0_conduit_end_CS_N,       //                               .CS_N
		output wire        cy7c67200_if_0_conduit_end_RST_N,      //                               .RST_N
		input  wire        cy7c67200_if_0_conduit_end_INT,        //                               .INT
		output wire        lcd_16207_0_external_RS,               //           lcd_16207_0_external.RS
		output wire        lcd_16207_0_external_RW,               //                               .RW
		inout  wire [7:0]  lcd_16207_0_external_data,             //                               .data
		output wire        lcd_16207_0_external_E,                //                               .E
		output wire [8:0]  led_green_external_connection_export,  //  led_green_external_connection.export
		output wire [17:0] led_red_external_connection_export,    //    led_red_external_connection.export
		output wire [12:0] sdram_0_wire_addr,                     //                   sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                       //                               .ba
		output wire        sdram_0_wire_cas_n,                    //                               .cas_n
		output wire        sdram_0_wire_cke,                      //                               .cke
		output wire        sdram_0_wire_cs_n,                     //                               .cs_n
		inout  wire [31:0] sdram_0_wire_dq,                       //                               .dq
		output wire [3:0]  sdram_0_wire_dqm,                      //                               .dqm
		output wire        sdram_0_wire_ras_n,                    //                               .ras_n
		output wire        sdram_0_wire_we_n,                     //                               .we_n
		output wire [6:0]  seg7_display_conduit_end_oSEG0,        //       seg7_display_conduit_end.oSEG0
		output wire [6:0]  seg7_display_conduit_end_oSEG1,        //                               .oSEG1
		output wire [6:0]  seg7_display_conduit_end_oSEG2,        //                               .oSEG2
		output wire [6:0]  seg7_display_conduit_end_oSEG3,        //                               .oSEG3
		output wire [6:0]  seg7_display_conduit_end_oSEG4,        //                               .oSEG4
		output wire [6:0]  seg7_display_conduit_end_oSEG5,        //                               .oSEG5
		output wire [6:0]  seg7_display_conduit_end_oSEG6,        //                               .oSEG6
		output wire [6:0]  seg7_display_conduit_end_oSEG7,        //                               .oSEG7
		input  wire [17:0] switch_pio_external_connection_export  // switch_pio_external_connection.export
	);

	wire  [31:0] cpu_0_data_master_readdata;                                    // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_waitrequest;                                 // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire         cpu_0_data_master_debugaccess;                                 // cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire  [27:0] cpu_0_data_master_address;                                     // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;                                  // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_0_data_master_read;                                        // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire         cpu_0_data_master_write;                                       // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                                   // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [31:0] cpu_0_instruction_master_readdata;                             // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [27:0] cpu_0_instruction_master_address;                              // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                                 // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire         cpu_0_instruction_master_readdatavalid;                        // mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;      // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;   // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_readdata;              // cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest;           // cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess;           // mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_0_debug_mem_slave_address;               // mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_read;                  // mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_0_debug_mem_slave_byteenable;            // mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_write;                 // mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_writedata;             // mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata;      // mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest;   // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid; // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire         mm_interconnect_0_sdram_0_s1_chipselect;                       // mm_interconnect_0:sdram_0_s1_chipselect -> sdram_0:az_cs
	wire  [31:0] mm_interconnect_0_sdram_0_s1_readdata;                         // sdram_0:za_data -> mm_interconnect_0:sdram_0_s1_readdata
	wire         mm_interconnect_0_sdram_0_s1_waitrequest;                      // sdram_0:za_waitrequest -> mm_interconnect_0:sdram_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_0_s1_address;                          // mm_interconnect_0:sdram_0_s1_address -> sdram_0:az_addr
	wire         mm_interconnect_0_sdram_0_s1_read;                             // mm_interconnect_0:sdram_0_s1_read -> sdram_0:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_0_s1_byteenable;                       // mm_interconnect_0:sdram_0_s1_byteenable -> sdram_0:az_be_n
	wire         mm_interconnect_0_sdram_0_s1_readdatavalid;                    // sdram_0:za_valid -> mm_interconnect_0:sdram_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_0_s1_write;                            // mm_interconnect_0:sdram_0_s1_write -> sdram_0:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_0_s1_writedata;                        // mm_interconnect_0:sdram_0_s1_writedata -> sdram_0:az_data
	wire         mm_clock_crossing_bridge_0_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_0_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire         mm_clock_crossing_bridge_0_m0_debugaccess;                     // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_0_m0_address;                         // mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_address
	wire         mm_clock_crossing_bridge_0_m0_read;                            // mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_read
	wire   [3:0] mm_clock_crossing_bridge_0_m0_byteenable;                      // mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_byteenable
	wire         mm_clock_crossing_bridge_0_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_0_m0_writedata;                       // mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_writedata
	wire         mm_clock_crossing_bridge_0_m0_write;                           // mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_write
	wire   [0:0] mm_clock_crossing_bridge_0_m0_burstcount;                      // mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_burstcount
	wire         mm_interconnect_1_seg7_display_avalon_slave_write;             // mm_interconnect_1:SEG7_Display_avalon_slave_write -> SEG7_Display:iWR
	wire  [31:0] mm_interconnect_1_seg7_display_avalon_slave_writedata;         // mm_interconnect_1:SEG7_Display_avalon_slave_writedata -> SEG7_Display:iDIG
	wire   [7:0] mm_interconnect_1_lcd_16207_0_control_slave_readdata;          // lcd_16207_0:readdata -> mm_interconnect_1:lcd_16207_0_control_slave_readdata
	wire   [1:0] mm_interconnect_1_lcd_16207_0_control_slave_address;           // mm_interconnect_1:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	wire         mm_interconnect_1_lcd_16207_0_control_slave_read;              // mm_interconnect_1:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	wire         mm_interconnect_1_lcd_16207_0_control_slave_begintransfer;     // mm_interconnect_1:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	wire         mm_interconnect_1_lcd_16207_0_control_slave_write;             // mm_interconnect_1:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	wire   [7:0] mm_interconnect_1_lcd_16207_0_control_slave_writedata;         // mm_interconnect_1:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	wire         mm_interconnect_1_cy7c67200_if_0_hpi_chipselect;               // mm_interconnect_1:CY7C67200_IF_0_hpi_chipselect -> CY7C67200_IF_0:iCS_N
	wire  [31:0] mm_interconnect_1_cy7c67200_if_0_hpi_readdata;                 // CY7C67200_IF_0:oDATA -> mm_interconnect_1:CY7C67200_IF_0_hpi_readdata
	wire   [1:0] mm_interconnect_1_cy7c67200_if_0_hpi_address;                  // mm_interconnect_1:CY7C67200_IF_0_hpi_address -> CY7C67200_IF_0:iADDR
	wire         mm_interconnect_1_cy7c67200_if_0_hpi_read;                     // mm_interconnect_1:CY7C67200_IF_0_hpi_read -> CY7C67200_IF_0:iRD_N
	wire         mm_interconnect_1_cy7c67200_if_0_hpi_write;                    // mm_interconnect_1:CY7C67200_IF_0_hpi_write -> CY7C67200_IF_0:iWR_N
	wire  [31:0] mm_interconnect_1_cy7c67200_if_0_hpi_writedata;                // mm_interconnect_1:CY7C67200_IF_0_hpi_writedata -> CY7C67200_IF_0:iDATA
	wire         mm_interconnect_1_timer_0_s1_chipselect;                       // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_1_timer_0_s1_readdata;                         // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_0_s1_address;                          // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_1_timer_0_s1_write;                            // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_1_timer_0_s1_writedata;                        // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_1_switch_pio_s1_readdata;                      // switch_pio:readdata -> mm_interconnect_1:switch_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_switch_pio_s1_address;                       // mm_interconnect_1:switch_pio_s1_address -> switch_pio:address
	wire         mm_interconnect_1_button_pio_s1_chipselect;                    // mm_interconnect_1:button_pio_s1_chipselect -> button_pio:chipselect
	wire  [31:0] mm_interconnect_1_button_pio_s1_readdata;                      // button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_button_pio_s1_address;                       // mm_interconnect_1:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_1_button_pio_s1_write;                         // mm_interconnect_1:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_1_button_pio_s1_writedata;                     // mm_interconnect_1:button_pio_s1_writedata -> button_pio:writedata
	wire         mm_interconnect_1_led_green_s1_chipselect;                     // mm_interconnect_1:led_green_s1_chipselect -> led_green:chipselect
	wire  [31:0] mm_interconnect_1_led_green_s1_readdata;                       // led_green:readdata -> mm_interconnect_1:led_green_s1_readdata
	wire   [1:0] mm_interconnect_1_led_green_s1_address;                        // mm_interconnect_1:led_green_s1_address -> led_green:address
	wire         mm_interconnect_1_led_green_s1_write;                          // mm_interconnect_1:led_green_s1_write -> led_green:write_n
	wire  [31:0] mm_interconnect_1_led_green_s1_writedata;                      // mm_interconnect_1:led_green_s1_writedata -> led_green:writedata
	wire         mm_interconnect_1_led_red_s1_chipselect;                       // mm_interconnect_1:led_red_s1_chipselect -> led_red:chipselect
	wire  [31:0] mm_interconnect_1_led_red_s1_readdata;                         // led_red:readdata -> mm_interconnect_1:led_red_s1_readdata
	wire   [1:0] mm_interconnect_1_led_red_s1_address;                          // mm_interconnect_1:led_red_s1_address -> led_red:address
	wire         mm_interconnect_1_led_red_s1_write;                            // mm_interconnect_1:led_red_s1_write -> led_red:write_n
	wire  [31:0] mm_interconnect_1_led_red_s1_writedata;                        // mm_interconnect_1:led_red_s1_writedata -> led_red:writedata
	wire         mm_interconnect_1_timer_1_s1_chipselect;                       // mm_interconnect_1:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_1_timer_1_s1_readdata;                         // timer_1:readdata -> mm_interconnect_1:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_1_s1_address;                          // mm_interconnect_1:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_1_timer_1_s1_write;                            // mm_interconnect_1:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_1_timer_1_s1_writedata;                        // mm_interconnect_1:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver1_irq;                                      // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_0_irq_irq;                                                 // irq_mapper:sender_irq -> cpu_0:irq
	wire         irq_mapper_receiver0_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                 // CY7C67200_IF_0:oINT -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                      // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                             // timer_0:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver3_irq;                                      // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                             // timer_1:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver4_irq;                                      // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                             // button_pio:irq -> irq_synchronizer_003:receiver_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [CY7C67200_IF_0:iRST_N, SEG7_Display:iRST_N, button_pio:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, lcd_16207_0:reset_n, led_green:reset_n, led_red:reset_n, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset, switch_pio:reset_n, timer_0:reset_n, timer_1:reset_n]
	wire         cpu_0_debug_reset_request_reset;                               // cpu_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [cpu_0:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, jtag_uart_0:rst_n, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                        // rst_controller_001:reset_req -> [cpu_0:reset_req, rst_translator:reset_req_in]

	CY7C67200_IF cy7c67200_if_0 (
		.oDATA     (mm_interconnect_1_cy7c67200_if_0_hpi_readdata),    //              hpi.readdata
		.iADDR     (mm_interconnect_1_cy7c67200_if_0_hpi_address),     //                 .address
		.iRD_N     (~mm_interconnect_1_cy7c67200_if_0_hpi_read),       //                 .read_n
		.iWR_N     (~mm_interconnect_1_cy7c67200_if_0_hpi_write),      //                 .write_n
		.iCS_N     (~mm_interconnect_1_cy7c67200_if_0_hpi_chipselect), //                 .chipselect_n
		.iDATA     (mm_interconnect_1_cy7c67200_if_0_hpi_writedata),   //                 .writedata
		.iCLK      (clk_io_clk_in_clk),                                //       clock_sink.clk
		.iRST_N    (~rst_controller_reset_out_reset),                  // clock_sink_reset.reset_n
		.oINT      (irq_synchronizer_receiver_irq),                    // interrupt_sender.irq
		.HPI_DATA  (cy7c67200_if_0_conduit_end_DATA),                  //      conduit_end.export
		.HPI_ADDR  (cy7c67200_if_0_conduit_end_ADDR),                  //                 .export
		.HPI_RD_N  (cy7c67200_if_0_conduit_end_RD_N),                  //                 .export
		.HPI_WR_N  (cy7c67200_if_0_conduit_end_WR_N),                  //                 .export
		.HPI_CS_N  (cy7c67200_if_0_conduit_end_CS_N),                  //                 .export
		.HPI_RST_N (cy7c67200_if_0_conduit_end_RST_N),                 //                 .export
		.HPI_INT   (cy7c67200_if_0_conduit_end_INT)                    //                 .export
	);

	SEG7_LUT_8 seg7_display (
		.iCLK   (clk_io_clk_in_clk),                                     //          clk.clk
		.iRST_N (~rst_controller_reset_out_reset),                       //    clk_reset.reset_n
		.iWR    (mm_interconnect_1_seg7_display_avalon_slave_write),     // avalon_slave.write
		.iDIG   (mm_interconnect_1_seg7_display_avalon_slave_writedata), //             .writedata
		.oSEG0  (seg7_display_conduit_end_oSEG0),                        //  conduit_end.export
		.oSEG1  (seg7_display_conduit_end_oSEG1),                        //             .export
		.oSEG2  (seg7_display_conduit_end_oSEG2),                        //             .export
		.oSEG3  (seg7_display_conduit_end_oSEG3),                        //             .export
		.oSEG4  (seg7_display_conduit_end_oSEG4),                        //             .export
		.oSEG5  (seg7_display_conduit_end_oSEG5),                        //             .export
		.oSEG6  (seg7_display_conduit_end_oSEG6),                        //             .export
		.oSEG7  (seg7_display_conduit_end_oSEG7)                         //             .export
	);

	DE2_115_Qsys_button_pio button_pio (
		.clk        (clk_io_clk_in_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_003_receiver_irq)           //                 irq.irq
	);

	DE2_115_Qsys_cpu_0 cpu_0 (
		.clk                                 (clk_100_clk_in_clk),                                  //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (cpu_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	DE2_115_Qsys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_100_clk_in_clk),                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	DE2_115_Qsys_lcd_16207_0 lcd_16207_0 (
		.reset_n       (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.clk           (clk_io_clk_in_clk),                                         //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_16207_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_16207_0_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_16207_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_16207_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_16207_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_16207_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_16207_0_external_RS),                                   //      external.export
		.LCD_RW        (lcd_16207_0_external_RW),                                   //              .export
		.LCD_data      (lcd_16207_0_external_data),                                 //              .export
		.LCD_E         (lcd_16207_0_external_E)                                     //              .export
	);

	DE2_115_Qsys_led_green led_green (
		.clk        (clk_io_clk_in_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_green_s1_readdata),   //                    .readdata
		.out_port   (led_green_external_connection_export)       // external_connection.export
	);

	DE2_115_Qsys_led_red led_red (
		.clk        (clk_io_clk_in_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_led_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_red_s1_readdata),   //                    .readdata
		.out_port   (led_red_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (clk_io_clk_in_clk),                                             //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                                // m0_reset.reset
		.s0_clk           (clk_100_clk_in_clk),                                            //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_Qsys_sdram_0 sdram_0 (
		.clk            (clk_100_clk_in_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),        // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                          //  wire.export
		.zs_ba          (sdram_0_wire_ba),                            //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                         //      .export
		.zs_cke         (sdram_0_wire_cke),                           //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                          //      .export
		.zs_dq          (sdram_0_wire_dq),                            //      .export
		.zs_dqm         (sdram_0_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_0_wire_we_n)                           //      .export
	);

	DE2_115_Qsys_switch_pio switch_pio (
		.clk      (clk_io_clk_in_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_switch_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_switch_pio_s1_readdata), //                    .readdata
		.in_port  (switch_pio_external_connection_export)     // external_connection.export
	);

	DE2_115_Qsys_timer_0 timer_0 (
		.clk        (clk_io_clk_in_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)        //   irq.irq
	);

	DE2_115_Qsys_timer_0 timer_1 (
		.clk        (clk_io_clk_in_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_1_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)        //   irq.irq
	);

	DE2_115_Qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_100_clk_clk                             (clk_100_clk_in_clk),                                            //                       clk_100_clk.clk
		.cpu_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                            // cpu_0_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                   (cpu_0_data_master_address),                                     //                 cpu_0_data_master.address
		.cpu_0_data_master_waitrequest               (cpu_0_data_master_waitrequest),                                 //                                  .waitrequest
		.cpu_0_data_master_byteenable                (cpu_0_data_master_byteenable),                                  //                                  .byteenable
		.cpu_0_data_master_read                      (cpu_0_data_master_read),                                        //                                  .read
		.cpu_0_data_master_readdata                  (cpu_0_data_master_readdata),                                    //                                  .readdata
		.cpu_0_data_master_write                     (cpu_0_data_master_write),                                       //                                  .write
		.cpu_0_data_master_writedata                 (cpu_0_data_master_writedata),                                   //                                  .writedata
		.cpu_0_data_master_debugaccess               (cpu_0_data_master_debugaccess),                                 //                                  .debugaccess
		.cpu_0_instruction_master_address            (cpu_0_instruction_master_address),                              //          cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest        (cpu_0_instruction_master_waitrequest),                          //                                  .waitrequest
		.cpu_0_instruction_master_read               (cpu_0_instruction_master_read),                                 //                                  .read
		.cpu_0_instruction_master_readdata           (cpu_0_instruction_master_readdata),                             //                                  .readdata
		.cpu_0_instruction_master_readdatavalid      (cpu_0_instruction_master_readdatavalid),                        //                                  .readdatavalid
		.cpu_0_debug_mem_slave_address               (mm_interconnect_0_cpu_0_debug_mem_slave_address),               //             cpu_0_debug_mem_slave.address
		.cpu_0_debug_mem_slave_write                 (mm_interconnect_0_cpu_0_debug_mem_slave_write),                 //                                  .write
		.cpu_0_debug_mem_slave_read                  (mm_interconnect_0_cpu_0_debug_mem_slave_read),                  //                                  .read
		.cpu_0_debug_mem_slave_readdata              (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),              //                                  .readdata
		.cpu_0_debug_mem_slave_writedata             (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),             //                                  .writedata
		.cpu_0_debug_mem_slave_byteenable            (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),            //                                  .byteenable
		.cpu_0_debug_mem_slave_waitrequest           (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest),           //                                  .waitrequest
		.cpu_0_debug_mem_slave_debugaccess           (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess),           //                                  .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),       //     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),         //                                  .write
		.jtag_uart_0_avalon_jtag_slave_read          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),          //                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),      //                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),     //                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),   //                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),    //                                  .chipselect
		.mm_clock_crossing_bridge_0_s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //     mm_clock_crossing_bridge_0_s0.address
		.mm_clock_crossing_bridge_0_s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //                                  .write
		.mm_clock_crossing_bridge_0_s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //                                  .read
		.mm_clock_crossing_bridge_0_s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //                                  .readdata
		.mm_clock_crossing_bridge_0_s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //                                  .writedata
		.mm_clock_crossing_bridge_0_s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //                                  .burstcount
		.mm_clock_crossing_bridge_0_s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //                                  .byteenable
		.mm_clock_crossing_bridge_0_s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //                                  .readdatavalid
		.mm_clock_crossing_bridge_0_s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //                                  .waitrequest
		.mm_clock_crossing_bridge_0_s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //                                  .debugaccess
		.sdram_0_s1_address                          (mm_interconnect_0_sdram_0_s1_address),                          //                        sdram_0_s1.address
		.sdram_0_s1_write                            (mm_interconnect_0_sdram_0_s1_write),                            //                                  .write
		.sdram_0_s1_read                             (mm_interconnect_0_sdram_0_s1_read),                             //                                  .read
		.sdram_0_s1_readdata                         (mm_interconnect_0_sdram_0_s1_readdata),                         //                                  .readdata
		.sdram_0_s1_writedata                        (mm_interconnect_0_sdram_0_s1_writedata),                        //                                  .writedata
		.sdram_0_s1_byteenable                       (mm_interconnect_0_sdram_0_s1_byteenable),                       //                                  .byteenable
		.sdram_0_s1_readdatavalid                    (mm_interconnect_0_sdram_0_s1_readdatavalid),                    //                                  .readdatavalid
		.sdram_0_s1_waitrequest                      (mm_interconnect_0_sdram_0_s1_waitrequest),                      //                                  .waitrequest
		.sdram_0_s1_chipselect                       (mm_interconnect_0_sdram_0_s1_chipselect)                        //                                  .chipselect
	);

	DE2_115_Qsys_mm_interconnect_1 mm_interconnect_1 (
		.clk_io_clk_clk                                                  (clk_io_clk_in_clk),                                         //                                                clk_io_clk.clk
		.mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_address                           (mm_clock_crossing_bridge_0_m0_address),                     //                             mm_clock_crossing_bridge_0_m0.address
		.mm_clock_crossing_bridge_0_m0_waitrequest                       (mm_clock_crossing_bridge_0_m0_waitrequest),                 //                                                          .waitrequest
		.mm_clock_crossing_bridge_0_m0_burstcount                        (mm_clock_crossing_bridge_0_m0_burstcount),                  //                                                          .burstcount
		.mm_clock_crossing_bridge_0_m0_byteenable                        (mm_clock_crossing_bridge_0_m0_byteenable),                  //                                                          .byteenable
		.mm_clock_crossing_bridge_0_m0_read                              (mm_clock_crossing_bridge_0_m0_read),                        //                                                          .read
		.mm_clock_crossing_bridge_0_m0_readdata                          (mm_clock_crossing_bridge_0_m0_readdata),                    //                                                          .readdata
		.mm_clock_crossing_bridge_0_m0_readdatavalid                     (mm_clock_crossing_bridge_0_m0_readdatavalid),               //                                                          .readdatavalid
		.mm_clock_crossing_bridge_0_m0_write                             (mm_clock_crossing_bridge_0_m0_write),                       //                                                          .write
		.mm_clock_crossing_bridge_0_m0_writedata                         (mm_clock_crossing_bridge_0_m0_writedata),                   //                                                          .writedata
		.mm_clock_crossing_bridge_0_m0_debugaccess                       (mm_clock_crossing_bridge_0_m0_debugaccess),                 //                                                          .debugaccess
		.button_pio_s1_address                                           (mm_interconnect_1_button_pio_s1_address),                   //                                             button_pio_s1.address
		.button_pio_s1_write                                             (mm_interconnect_1_button_pio_s1_write),                     //                                                          .write
		.button_pio_s1_readdata                                          (mm_interconnect_1_button_pio_s1_readdata),                  //                                                          .readdata
		.button_pio_s1_writedata                                         (mm_interconnect_1_button_pio_s1_writedata),                 //                                                          .writedata
		.button_pio_s1_chipselect                                        (mm_interconnect_1_button_pio_s1_chipselect),                //                                                          .chipselect
		.CY7C67200_IF_0_hpi_address                                      (mm_interconnect_1_cy7c67200_if_0_hpi_address),              //                                        CY7C67200_IF_0_hpi.address
		.CY7C67200_IF_0_hpi_write                                        (mm_interconnect_1_cy7c67200_if_0_hpi_write),                //                                                          .write
		.CY7C67200_IF_0_hpi_read                                         (mm_interconnect_1_cy7c67200_if_0_hpi_read),                 //                                                          .read
		.CY7C67200_IF_0_hpi_readdata                                     (mm_interconnect_1_cy7c67200_if_0_hpi_readdata),             //                                                          .readdata
		.CY7C67200_IF_0_hpi_writedata                                    (mm_interconnect_1_cy7c67200_if_0_hpi_writedata),            //                                                          .writedata
		.CY7C67200_IF_0_hpi_chipselect                                   (mm_interconnect_1_cy7c67200_if_0_hpi_chipselect),           //                                                          .chipselect
		.lcd_16207_0_control_slave_address                               (mm_interconnect_1_lcd_16207_0_control_slave_address),       //                                 lcd_16207_0_control_slave.address
		.lcd_16207_0_control_slave_write                                 (mm_interconnect_1_lcd_16207_0_control_slave_write),         //                                                          .write
		.lcd_16207_0_control_slave_read                                  (mm_interconnect_1_lcd_16207_0_control_slave_read),          //                                                          .read
		.lcd_16207_0_control_slave_readdata                              (mm_interconnect_1_lcd_16207_0_control_slave_readdata),      //                                                          .readdata
		.lcd_16207_0_control_slave_writedata                             (mm_interconnect_1_lcd_16207_0_control_slave_writedata),     //                                                          .writedata
		.lcd_16207_0_control_slave_begintransfer                         (mm_interconnect_1_lcd_16207_0_control_slave_begintransfer), //                                                          .begintransfer
		.led_green_s1_address                                            (mm_interconnect_1_led_green_s1_address),                    //                                              led_green_s1.address
		.led_green_s1_write                                              (mm_interconnect_1_led_green_s1_write),                      //                                                          .write
		.led_green_s1_readdata                                           (mm_interconnect_1_led_green_s1_readdata),                   //                                                          .readdata
		.led_green_s1_writedata                                          (mm_interconnect_1_led_green_s1_writedata),                  //                                                          .writedata
		.led_green_s1_chipselect                                         (mm_interconnect_1_led_green_s1_chipselect),                 //                                                          .chipselect
		.led_red_s1_address                                              (mm_interconnect_1_led_red_s1_address),                      //                                                led_red_s1.address
		.led_red_s1_write                                                (mm_interconnect_1_led_red_s1_write),                        //                                                          .write
		.led_red_s1_readdata                                             (mm_interconnect_1_led_red_s1_readdata),                     //                                                          .readdata
		.led_red_s1_writedata                                            (mm_interconnect_1_led_red_s1_writedata),                    //                                                          .writedata
		.led_red_s1_chipselect                                           (mm_interconnect_1_led_red_s1_chipselect),                   //                                                          .chipselect
		.SEG7_Display_avalon_slave_write                                 (mm_interconnect_1_seg7_display_avalon_slave_write),         //                                 SEG7_Display_avalon_slave.write
		.SEG7_Display_avalon_slave_writedata                             (mm_interconnect_1_seg7_display_avalon_slave_writedata),     //                                                          .writedata
		.switch_pio_s1_address                                           (mm_interconnect_1_switch_pio_s1_address),                   //                                             switch_pio_s1.address
		.switch_pio_s1_readdata                                          (mm_interconnect_1_switch_pio_s1_readdata),                  //                                                          .readdata
		.timer_0_s1_address                                              (mm_interconnect_1_timer_0_s1_address),                      //                                                timer_0_s1.address
		.timer_0_s1_write                                                (mm_interconnect_1_timer_0_s1_write),                        //                                                          .write
		.timer_0_s1_readdata                                             (mm_interconnect_1_timer_0_s1_readdata),                     //                                                          .readdata
		.timer_0_s1_writedata                                            (mm_interconnect_1_timer_0_s1_writedata),                    //                                                          .writedata
		.timer_0_s1_chipselect                                           (mm_interconnect_1_timer_0_s1_chipselect),                   //                                                          .chipselect
		.timer_1_s1_address                                              (mm_interconnect_1_timer_1_s1_address),                      //                                                timer_1_s1.address
		.timer_1_s1_write                                                (mm_interconnect_1_timer_1_s1_write),                        //                                                          .write
		.timer_1_s1_readdata                                             (mm_interconnect_1_timer_1_s1_readdata),                     //                                                          .readdata
		.timer_1_s1_writedata                                            (mm_interconnect_1_timer_1_s1_writedata),                    //                                                          .writedata
		.timer_1_s1_chipselect                                           (mm_interconnect_1_timer_1_s1_chipselect)                    //                                                          .chipselect
	);

	DE2_115_Qsys_irq_mapper irq_mapper (
		.clk           (clk_100_clk_in_clk),                 //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_0_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_io_clk_in_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_100_clk_in_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_io_clk_in_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_100_clk_in_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_io_clk_in_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_100_clk_in_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_io_clk_in_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_100_clk_in_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_100_clk_in_reset_reset_n),   // reset_in0.reset
		.reset_in1      (cpu_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_io_clk_in_clk),               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                // (terminated)
		.reset_req_in0  (1'b0),                            // (terminated)
		.reset_req_in1  (1'b0),                            // (terminated)
		.reset_in2      (1'b0),                            // (terminated)
		.reset_req_in2  (1'b0),                            // (terminated)
		.reset_in3      (1'b0),                            // (terminated)
		.reset_req_in3  (1'b0),                            // (terminated)
		.reset_in4      (1'b0),                            // (terminated)
		.reset_req_in4  (1'b0),                            // (terminated)
		.reset_in5      (1'b0),                            // (terminated)
		.reset_req_in5  (1'b0),                            // (terminated)
		.reset_in6      (1'b0),                            // (terminated)
		.reset_req_in6  (1'b0),                            // (terminated)
		.reset_in7      (1'b0),                            // (terminated)
		.reset_req_in7  (1'b0),                            // (terminated)
		.reset_in8      (1'b0),                            // (terminated)
		.reset_req_in8  (1'b0),                            // (terminated)
		.reset_in9      (1'b0),                            // (terminated)
		.reset_req_in9  (1'b0),                            // (terminated)
		.reset_in10     (1'b0),                            // (terminated)
		.reset_req_in10 (1'b0),                            // (terminated)
		.reset_in11     (1'b0),                            // (terminated)
		.reset_req_in11 (1'b0),                            // (terminated)
		.reset_in12     (1'b0),                            // (terminated)
		.reset_req_in12 (1'b0),                            // (terminated)
		.reset_in13     (1'b0),                            // (terminated)
		.reset_req_in13 (1'b0),                            // (terminated)
		.reset_in14     (1'b0),                            // (terminated)
		.reset_req_in14 (1'b0),                            // (terminated)
		.reset_in15     (1'b0),                            // (terminated)
		.reset_req_in15 (1'b0)                             // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clk_100_clk_in_reset_reset_n),          // reset_in0.reset
		.reset_in1      (cpu_0_debug_reset_request_reset),        // reset_in1.reset
		.clk            (clk_100_clk_in_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
