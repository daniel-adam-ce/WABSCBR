module sboxinst1(
	input [7:0] unboxed,
	output reg[7:0] boxed);
	
	always@(*) begin 
	case (unboxed)
	8'h00: boxed=8'h63;
	8'h01: boxed=8'h7c;
	8'h02: boxed=8'h77;
	8'h03: boxed=8'h7b;
	8'h04: boxed=8'hf2;
	8'h05: boxed=8'h6b;
	8'h06: boxed=8'h6f;
	8'h07: boxed=8'hc5;
	8'h08: boxed=8'h30;
	8'h09: boxed=8'h01;
	8'h0a: boxed=8'h67;
	8'h0b: boxed=8'h2b;
	8'h0c: boxed=8'hfe;
	8'h0d: boxed=8'hd7;
	8'h0e: boxed=8'hab;
	8'h0f: boxed=8'h76;
	8'h10: boxed=8'hca;
	8'h11: boxed=8'h82;
	8'h12: boxed=8'hc9;
	8'h13: boxed=8'h7d;
	8'h14: boxed=8'hfa;
	8'h15: boxed=8'h59;
	8'h16: boxed=8'h47;
	8'h17: boxed=8'hf0;
	8'h18: boxed=8'had;
	8'h19: boxed=8'hd4;
	8'h1a: boxed=8'ha2;
	8'h1b: boxed=8'haf;
	8'h1c: boxed=8'h9c;
	8'h1d: boxed=8'ha4;
	8'h1e: boxed=8'h72;
	8'h1f: boxed=8'hc0;
	8'h20: boxed=8'hb7;
	8'h21: boxed=8'hfd;
	8'h22: boxed=8'h93;
	8'h23: boxed=8'h26;
	8'h24: boxed=8'h36;
	8'h25: boxed=8'h3f;
	8'h26: boxed=8'hf7;
	8'h27: boxed=8'hcc;
	8'h28: boxed=8'h34;
	8'h29: boxed=8'ha5;
	8'h2a: boxed=8'he5;
	8'h2b: boxed=8'hf1;
	8'h2c: boxed=8'h71;
	8'h2d: boxed=8'hd8;
	8'h2e: boxed=8'h31;
	8'h2f: boxed=8'h15;
	8'h30: boxed=8'h04;
	8'h31: boxed=8'hc7;
	8'h32: boxed=8'h23;
	8'h33: boxed=8'hc3;
	8'h34: boxed=8'h18;
	8'h35: boxed=8'h96;
	8'h36: boxed=8'h05;
	8'h37: boxed=8'h9a;
	8'h38: boxed=8'h07;
	8'h39: boxed=8'h12;
	8'h3a: boxed=8'h80;
	8'h3b: boxed=8'he2;
	8'h3c: boxed=8'heb;
	8'h3d: boxed=8'h27;
	8'h3e: boxed=8'hb2;
	8'h3f: boxed=8'h75;
	8'h40: boxed=8'h09;
	8'h41: boxed=8'h83;
	8'h42: boxed=8'h2c;
	8'h43: boxed=8'h1a;
	8'h44: boxed=8'h1b;
	8'h45: boxed=8'h6e;
	8'h46: boxed=8'h5a;
	8'h47: boxed=8'ha0;
	8'h48: boxed=8'h52;
	8'h49: boxed=8'h3b;
	8'h4a: boxed=8'hd6;
	8'h4b: boxed=8'hb3;
	8'h4c: boxed=8'h29;
	8'h4d: boxed=8'he3;
	8'h4e: boxed=8'h2f;
	8'h4f: boxed=8'h84;
	8'h50: boxed=8'h53;
	8'h51: boxed=8'hd1;
	8'h52: boxed=8'h00;
	8'h53: boxed=8'hed;
	8'h54: boxed=8'h20;
	8'h55: boxed=8'hfc;
	8'h56: boxed=8'hb1;
	8'h57: boxed=8'h5b;
	8'h58: boxed=8'h6a;
	8'h59: boxed=8'hcb;
	8'h5a: boxed=8'hbe;
	8'h5b: boxed=8'h39;
	8'h5c: boxed=8'h4a;
	8'h5d: boxed=8'h4c;
	8'h5e: boxed=8'h58;
	8'h5f: boxed=8'hcf;
	8'h60: boxed=8'hd0;
	8'h61: boxed=8'hef;
	8'h62: boxed=8'haa;
	8'h63: boxed=8'hfb;
	8'h64: boxed=8'h43;
	8'h65: boxed=8'h4d;
	8'h66: boxed=8'h33;
	8'h67: boxed=8'h85;
	8'h68: boxed=8'h45;
	8'h69: boxed=8'hf9;
	8'h6a: boxed=8'h02;
	8'h6b: boxed=8'h7f;
	8'h6c: boxed=8'h50;
	8'h6d: boxed=8'h3c;
	8'h6e: boxed=8'h9f;
	8'h6f: boxed=8'ha8;
	8'h70: boxed=8'h51;
	8'h71: boxed=8'ha3;
	8'h72: boxed=8'h40;
	8'h73: boxed=8'h8f;
	8'h74: boxed=8'h92;
	8'h75: boxed=8'h9d;
	8'h76: boxed=8'h38;
	8'h77: boxed=8'hf5;
	8'h78: boxed=8'hbc;
	8'h79: boxed=8'hb6;
	8'h7a: boxed=8'hda;
	8'h7b: boxed=8'h21;
	8'h7c: boxed=8'h10;
	8'h7d: boxed=8'hff;
	8'h7e: boxed=8'hf3;
	8'h7f: boxed=8'hd2;
	8'h80: boxed=8'hcd;
	8'h81: boxed=8'h0c;
	8'h82: boxed=8'h13;
	8'h83: boxed=8'hec;
	8'h84: boxed=8'h5f;
	8'h85: boxed=8'h97;
	8'h86: boxed=8'h44;
	8'h87: boxed=8'h17;
	8'h88: boxed=8'hc4;
	8'h89: boxed=8'ha7;
	8'h8a: boxed=8'h7e;
	8'h8b: boxed=8'h3d;
	8'h8c: boxed=8'h64;
	8'h8d: boxed=8'h5d;
	8'h8e: boxed=8'h19;
	8'h8f: boxed=8'h73;
	8'h90: boxed=8'h60;
	8'h91: boxed=8'h81;
	8'h92: boxed=8'h4f;
	8'h93: boxed=8'hdc;
	8'h94: boxed=8'h22;
	8'h95: boxed=8'h2a;
	8'h96: boxed=8'h90;
	8'h97: boxed=8'h88;
	8'h98: boxed=8'h46;
	8'h99: boxed=8'hee;
	8'h9a: boxed=8'hb8;
	8'h9b: boxed=8'h14;
	8'h9c: boxed=8'hde;
	8'h9d: boxed=8'h5e;
	8'h9e: boxed=8'h0b;
	8'h9f: boxed=8'hdb;
	8'ha0: boxed=8'he0;
	8'ha1: boxed=8'h32;
	8'ha2: boxed=8'h3a;
	8'ha3: boxed=8'h0a;
	8'ha4: boxed=8'h49;
	8'ha5: boxed=8'h06;
	8'ha6: boxed=8'h24;
	8'ha7: boxed=8'h5c;
	8'ha8: boxed=8'hc2;
	8'ha9: boxed=8'hd3;
	8'haa: boxed=8'hac;
	8'hab: boxed=8'h62;
	8'hac: boxed=8'h91;
	8'had: boxed=8'h95;
	8'hae: boxed=8'he4;
	8'haf: boxed=8'h79;
	8'hb0: boxed=8'he7;
	8'hb1: boxed=8'hc8;
	8'hb2: boxed=8'h37;
	8'hb3: boxed=8'h6d;
	8'hb4: boxed=8'h8d;
	8'hb5: boxed=8'hd5;
	8'hb6: boxed=8'h4e;
	8'hb7: boxed=8'ha9;
	8'hb8: boxed=8'h6c;
	8'hb9: boxed=8'h56;
	8'hba: boxed=8'hf4;
	8'hbb: boxed=8'hea;
	8'hbc: boxed=8'h65;
	8'hbd: boxed=8'h7a;
	8'hbe: boxed=8'hae;
	8'hbf: boxed=8'h08;
	8'hc0: boxed=8'hba;
	8'hc1: boxed=8'h78;
	8'hc2: boxed=8'h25;
	8'hc3: boxed=8'h2e;
	8'hc4: boxed=8'h1c;
	8'hc5: boxed=8'ha6;
	8'hc6: boxed=8'hb4;
	8'hc7: boxed=8'hc6;
	8'hc8: boxed=8'he8;
	8'hc9: boxed=8'hdd;
	8'hca: boxed=8'h74;
	8'hcb: boxed=8'h1f;
	8'hcc: boxed=8'h4b;
	8'hcd: boxed=8'hbd;
	8'hce: boxed=8'h8b;
	8'hcf: boxed=8'h8a;
	8'hd0: boxed=8'h70;
	8'hd1: boxed=8'h3e;
	8'hd2: boxed=8'hb5;
	8'hd3: boxed=8'h66;
	8'hd4: boxed=8'h48;
	8'hd5: boxed=8'h03;
	8'hd6: boxed=8'hf6;
	8'hd7: boxed=8'h0e;
	8'hd8: boxed=8'h61;
	8'hd9: boxed=8'h35;
	8'hda: boxed=8'h57;
	8'hdb: boxed=8'hb9;
	8'hdc: boxed=8'h86;
	8'hdd: boxed=8'hc1;
	8'hde: boxed=8'h1d;
	8'hdf: boxed=8'h9e;
	8'he0: boxed=8'he1;
	8'he1: boxed=8'hf8;
	8'he2: boxed=8'h98;
	8'he3: boxed=8'h11;
	8'he4: boxed=8'h69;
	8'he5: boxed=8'hd9;
	8'he6: boxed=8'h8e;
	8'he7: boxed=8'h94;
	8'he8: boxed=8'h9b;
	8'he9: boxed=8'h1e;
	8'hea: boxed=8'h87;
	8'heb: boxed=8'he9;
	8'hec: boxed=8'hce;
	8'hed: boxed=8'h55;
	8'hee: boxed=8'h28;
	8'hef: boxed=8'hdf;
	8'hf0: boxed=8'h8c;
	8'hf1: boxed=8'ha1;
	8'hf2: boxed=8'h89;
	8'hf3: boxed=8'h0d;
	8'hf4: boxed=8'hbf;
	8'hf5: boxed=8'he6;
	8'hf6: boxed=8'h42;
	8'hf7: boxed=8'h68;
	8'hf8: boxed=8'h41;
	8'hf9: boxed=8'h99;
	8'hfa: boxed=8'h2d;
	8'hfb: boxed=8'h0f;
	8'hfc: boxed=8'hb0;
	8'hfd: boxed=8'h54;
	8'hfe: boxed=8'hbb;
	8'hff: boxed=8'h16;


	endcase
end
endmodule 
